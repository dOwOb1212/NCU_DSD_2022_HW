module D2_top(hsync, vsync, vga_r, vga_g, vga_b, LedOut, L_SevenSegOut, R_SevenSegOut, Enable, key_clk, key_data, S2, clk, reset, pclk);
output  hsync,vsync;
output  [7:0] Enable;
output  [3:0] vga_r, vga_g, vga_b;
output  [15:0] LedOut;
output  [6:0] L_SevenSegOut, R_SevenSegOut;
input   clk, reset, S2, key_clk, key_data, pclk;
wire f_clk, Led_clk, i_clk, snake_clk, SevenSeg_clk, c_clk, touchEdge, touchSelf, touchPoison, Touch_I_Fruit, Touch_N_Fruit, fruit, Long_enough, Touchbarrier;
wire [3:0] poison_x, poison_y, I_fruit_x, I_fruit_y, N_fruit_x, N_fruit_y;
wire [39:0] snake_x, snake_y; 
wire [2:0] NS, countDown;
wire [3:0] score100, score10, score1;
wire [1:0] direct;
wire [3:0] enable;
wire up, down, left, right, Q, start, key_state;
assign Enable = {enable,enable};
clkDivider u0(f_clk, Led_clk, i_clk, snake_clk, c_clk, SevenSeg_clk, clk, reset);
state u1 (NS, reset, clk, start, Long_enough, touchEdge, touchPoison, touchSelf, Touch_I_Fruit, Touchbarrier, countDown);
TouchPoison u3(touchPoison, snake_x[39:36], snake_y[39:36], NS, poison_x, poison_y);
TouchSelf u4(touchSelf, snake_x, snake_y);
TouchFruit u5(Touch_N_Fruit, Touch_I_Fruit, N_fruit_x, I_fruit_x, I_fruit_y, N_fruit_y, snake_x[39:36], snake_y[39:36]);
SnakeMove u6(flag, touchEdge, direct, snake_x, snake_y, NS, up, down, left, right, N_fruit_x, N_fruit_y, snake_clk, clk, reset, key_state);
I_fruit u7(I_fruit_x, I_fruit_y, NS, snake_x, snake_y, poison_x, poison_y, N_fruit_x, N_fruit_y, Q, Touch_I_fruit, clk, f_clk, reset, key_state);
N_fruit u8(fruit, N_fruit_x, N_fruit_y, I_fruit_x, I_fruit_y, Touch_N_Fruit, snake_x, snake_y, poison_x, poison_y, clk, f_clk, reset);
poison u9(poison_x, poison_y, NS, touchPoison, clk, reset);
VGA_display u10(pclk, clk, reset, start, hsync, vsync, vga_r, vga_g, vga_b, N_fruit_x, N_fruit_y, fruit, snake_y, snake_x, I_fruit_x, I_fruit_y, poison_x, poison_y, NS, flag);
CountDown u11(countDown, NS, c_clk, reset);
Score u12(score100, score10, score1, Touch_N_Fruit, NS, clk, reset);
SevenSegShow u13(L_SevenSegOut, R_SevenSegOut, enable, countDown, score100, score10, score1, NS, SevenSeg_clk, reset);
LedShow u14(LedOut, NS, Led_clk, reset);
Size u15(Long_enough, snake_x, snake_y);
TouchBarrier u16(Touchbarrier, snake_x[39:36], snake_y[39:36]);
keyboard u17(clk,reset,key_clk,key_data,up, left,down,right,Q,key_state);
debounce_D2 u18(S2, clk,reset, start);
endmodule
