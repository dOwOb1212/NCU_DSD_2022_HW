module Top(goRight, goLeft, clk, reset, start);
input goRight, goLeft, clk, reset, start;
wire [1:0]state;
wire OnElevator, OnElevator1, OnElevator2, OnElevator3, touch, drop, clk, reset, Key, goal;
wire [1:0]Chance;
wire [3:0]E1_yloc;
wire [3:0]E2_yloc;
wire [3:0]E3_yloc;
wire [3:0]E1_Yinit = 4'b0010;
wire [3:0]E2_Yinit = 4'b0110;
wire [3:0]E3_Yinit = 4'b1010;
wire [3:0]N_xloc;
wire [3:0]N_yloc;
wire [3:0]S1_yloc; 
wire [3:0]S2_yloc; 
wire [3:0]S3_yloc;
wire [3:0]S1_Yinit = 4'b1000;
wire [3:0]S2_Yinit = 4'b0101;
wire [3:0]S3_Yinit = 4'b0010;
wire [6:0]Score;
State State(state[1:0], N_xloc[3:0], N_yloc[3:0], Chance[1:0], start, OnElevator, touch, drop, clk, reset, goRight, goLeft);
Elevator Elevator1(E1_yloc[3:0], E1_Yinit[3:0], clk, reset, start);
Elevator Elevator2(E2_yloc[3:0], E2_Yinit[3:0], clk, reset, start);
Elevator Elevator3(E3_yloc[3:0], E3_Yinit[3:0], clk, reset, start);
OnElevation OnElevation1(OnElevator1, N_xloc[3:0], N_yloc[3:0], E1_yloc[3:0], goRight, goLeft);
OnElevation OnElevation2(OnElevator2, N_xloc[3:0], N_yloc[3:0], E2_yloc[3:0], goRight, goLeft);
OnElevation OnElevation3(OnElevator3, N_xloc[3:0], N_yloc[3:0], E3_yloc[3:0], goRight, goLeft);
Shuriken Shuriken1(S1_yloc[3:0], S1_Yinit[3:0], clk, reset);
Shuriken Shuriken2(S2_yloc[3:0], S2_Yinit[3:0], clk, reset);
Shuriken Shuriken3(S3_yloc[3:0], S3_Yinit[3:0], clk, reset);
Touch Touch(touch, N_xloc[3:0], N_yloc[3:0], S1_yloc[3:0], S2_yloc[3:0], S3_yloc[3:0]);
Drop Drop(drop, N_xloc[3:0], N_yloc[3:0], goRight, goLeft, E1_yloc[3:0], E2_yloc[3:0], E3_yloc[3:0]);
key key(Key, N_xloc[3:0], N_yloc[3:0]);
Goal Goal(goal, N_xloc[3:0], N_yloc[3:0]);
score score(Score[6:0], Key, goal);
assign OnElevator = OnElevator1 | OnElevator2 | OnElevator3;
endmodule
